--Johnny Li
--EEL4712 Digital Design
--Lab 7: top_level

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity top_level is
    port (
        clk50MHz : in  std_logic;
        switch   : in  std_logic_vector(9 downto 0);
        button   : in  std_logic_vector(1 downto 0);
        led0     : out std_logic_vector(6 downto 0);
        led0_dp  : out std_logic;
        led1     : out std_logic_vector(6 downto 0);
        led1_dp  : out std_logic;
        led2     : out std_logic_vector(6 downto 0);
        led2_dp  : out std_logic;
        led3     : out std_logic_vector(6 downto 0);
        led3_dp  : out std_logic;
        led4     : out std_logic_vector(6 downto 0);
        led4_dp  : out std_logic;
        led5     : out std_logic_vector(6 downto 0);
        led5_dp  : out std_logic
        );
end top_level;

architecture STR of top_level is

component decoder7seg
	port (
		input  : in  std_logic_vector(3 downto 0);
		output : out std_logic_vector(6 downto 0));
end component;

constant C0 : std_logic_vector(3 downto 0) := (others => '0');

signal outport0,intemp	: std_logic_vector(31 downto 0);
signal b0, in0, in1 : std_logic;
signal temp : std_logic_vector(31 downto 9);

begin  -- STR

	--b0 <= button(0);	--GCD
	b0 <= not button(0);	--bubble_sort
	in0 <= not switch(9) and not button(1);
	in1 <= switch(9) and not button(1);
	temp <= (others => '0');
	intemp <= temp & switch(8 downto 0);
    U_MIPS : entity work.mips
	port map (
		clk	=> clk50MHz,
		rst	=> b0,	
		Inport0_en => in0,
		Inport1_en => in1,
		InPort => intemp,
		OutPort	=> OutPort0
		);

    U_LED5 : decoder7seg port map (
        input  => C0,
        output => led5);

    U_LED4 : decoder7seg port map (
        input  => C0,
        output => led4);
    
    U_LED3 : decoder7seg port map (
        input  => OutPort0(15 downto 12),
        output => led3);

    U_LED2 : decoder7seg port map (
        input  => OutPort0(11 downto 8),
        output => led2);
    
    U_LED1 : decoder7seg port map (
        input  => OutPort0(7 downto 4),
        output => led1);

    U_LED0 : decoder7seg port map (
        input  => OutPort0(3 downto 0),
        output => led0);
    
    led5_dp <= '1';
    led4_dp <= '1';
    led3_dp <= '1';
    led2_dp <= '1';
    led1_dp <= '1';
    led0_dp <= '1';

end STR;